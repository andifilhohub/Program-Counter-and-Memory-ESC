`include "gram4k.v"

module tb_gram4k;
    // Relógio
    reg relogio_tb;
    
    // Sinal de habilitação
    reg habilita_tb;
    
    // Entradas e saída
    reg [15:0] dado_tb;
    reg [11:0] endereco_tb;  // 12 bits para endereçamento de 4k palavras
    wire [15:0] resultado_tb;

    // Unidade sob teste
    minha_ram4k instancia_ram (
        .dado_in(dado_tb),
        .endereco_in(endereco_tb),
        .habilita_in(habilita_tb),
        .relogio_in(relogio_tb),
        .dado_out(resultado_tb)
    );

    initial begin
        $display("Simulação personalizada da RAM 4K");
        $dumpfile("signals.vcd");
        $dumpvars(0, tb_gram4k);

        // Inicialização
        relogio_tb = 0;
        habilita_tb = 0;
        dado_tb = 16'b0000000000000000;
        endereco_tb = 12'b000000000000;
        
        // Teste escrevendo em diferentes endereços
        #1  habilita_tb = 1; dado_tb = 16'b1010101010101010; endereco_tb = 12'd0;
        #2  habilita_tb = 1; dado_tb = 16'b0101010101010101; endereco_tb = 12'd1;
        #2  habilita_tb = 1; dado_tb = 16'b1111000011110000; endereco_tb = 12'd2;
        #2  habilita_tb = 1; dado_tb = 16'b0000111100001111; endereco_tb = 12'd3;
        #2  habilita_tb = 1; dado_tb = 16'b1111111100000000; endereco_tb = 12'd4;
        #2  habilita_tb = 1; dado_tb = 16'b0000000011111111; endereco_tb = 12'd5;
        #2  habilita_tb = 1; dado_tb = 16'b1010101001010101; endereco_tb = 12'd100;
        #2  habilita_tb = 1; dado_tb = 16'b0101010110101010; endereco_tb = 12'd200;
        #2  habilita_tb = 1; dado_tb = 16'b1100110011001100; endereco_tb = 12'd300; 
        #2  habilita_tb = 1; dado_tb = 16'b0011001100110011; endereco_tb = 12'd400; 
        #2  habilita_tb = 1; dado_tb = 16'b1010010110100101; endereco_tb = 12'd500; 
        #2  habilita_tb = 1; dado_tb = 16'b0101101001011010; endereco_tb = 12'd4095; 

        // Teste de leitura dos registradores
        #2  habilita_tb = 0; endereco_tb = 12'd0;
        #2  endereco_tb = 12'd1; 
        #2  endereco_tb = 12'd2; 
        #2  endereco_tb = 12'd3; 
        #2  endereco_tb = 12'd4; 
        #2  endereco_tb = 12'd5; 
        #2  endereco_tb = 12'd100; 
        #2  endereco_tb = 12'd200; 
        #2  endereco_tb = 12'd300; 
        #2  endereco_tb = 12'd400; 
        #2  endereco_tb = 12'd500; 
        #2  endereco_tb = 12'd4095; 

        // Teste de atualização com habilita=0
        #2  habilita_tb = 0; dado_tb = 16'b1111111111111111; endereco_tb = 12'd0; // Não deve alterar
        #2  endereco_tb = 12'd0; // Verifica se o valor não foi alterado

        // Teste de atualização com habilita=1
        #2  habilita_tb = 1; dado_tb = 16'b1111111111111111; endereco_tb = 12'd0; // Deve alterar
        #2  habilita_tb = 0; endereco_tb = 12'd0; // Verifica a alteração

        #5  $finish;
    end

    initial begin
        $monitor("Tempo: %0t | Habilita: %b | Endereco: %3d | Dado: %b | Resultado: %b", $time, habilita_tb, endereco_tb, dado_tb, resultado_tb);
    end

    always #1 relogio_tb = ~relogio_tb;
    
endmodule